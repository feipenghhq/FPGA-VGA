../vga_core/vga_timing.svh